var SHUTDOWN = "Stäng av?",
OK = "OK",
CANCEL = "Avbryt",
CONFIGURATION = "Konfiguration",
UPLOAD_ERROR_FILETYPE = "Filen är inte tillåtet bildformat",
UPLOAD_ERROR_FILESIZE = "Maximalt tillåten storlek är 2MB";

